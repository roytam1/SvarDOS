#
# This is a localization file for the SvarDOS INSTALL program
# Detta �r en localiseringsfil f�r SvarDOSs INSTALLprogram
#
# Language..: Swedish
# Translator: Martin Str�mberg
#

### COMMON STUFF: TITLE BAR AND MULTIPLE CHOICE STRINGS ###
### GEMENSAMMA SAKER: TITLE-BAR AND MULTIPLA-VALSTR�NGAR ###
#0.0:SVARDOS INSTALLATION
0.0:SVARDOS INSTALLATION
#0.1:Install SvarDOS
0.1:Installera SvarDOS
#0.2:Quit to DOS
0.2:Avsluta till DOS
#0.3:Create a partition automatically
0.3:Skapa en partition automatiskt
#0.4:Run the FDISK partitioning tool
0.4:K�r FDISK-partitioneringsverktyget
#0.5:Press any key...
0.5:Tryck p� en tangent...
# Every string below must be at most 78 characters long! (used in status bar)
# Varje str�ng nedan m�ste vara som mest 78 bokst�ver l�ng (anv�nds i statusbaren)
#0.10:Up/Down = Select entry | Enter = Confirm choice | ESC = Previous screen
0.10:Upp/Ner = V�lj rad | Enter = Bekr�fta val | ESC = F�reg�ende sk�rm
#0.11:Up/Down = Select entry | Enter = Confirm choice | ESC = Quit to DOS
0.11:Up/Down = V�lj rad | Enter = Bekr�fta val | ESC = Avsluta till DOS

### LANGUAGE SELECTION & KEYBOARD LAYOUT SCREENS ###
### SPR�KVAL & TANGENTBORDSLAYOUTSK�RMAR ###
#1.0:Welcome to SvarDOS
1.0:V�lkommen till SvarDOS
#1.1:Please select your preferred language from the list below:
1.1:V�nligen v�lj spr�ket du vill anv�nda fr�n listan nedan:
#1.5:SvarDOS supports different keyboard layouts. Choose the keyboard layout that you want.
1.5:SvarDOS st�djer olika tangentbordslayouter. V�lj tangentbordslayouten som du vill ha.

### WELCOME SCREEN ###
### V�LKOMSTSK�RM ###
#2.0:You are about to install SvarDOS: a free, MS-DOS compatible operating system based on FreeDOS. SvarDOS comes with a variety of third-party applications.\n\nWARNING: If your PC has another operating system installed, this other system might be unable to boot once SvarDOS is installed.
2.0:Du ska just till att installera SvarDOS: ett fritt, MS-DOS-kompatibelt operativsystem baserat p� FreeDOS. SvarDOS kommer med en samling olika tredjepartsapplikationer.\n\nVARNING: Om din PC har ett annat operativsystem intstallerat, kanske detta andra system inte kan boota n�r v�l SvarDOS har installerats.

### DISK SETUP ###
### DISKSETUP ###
#3.0:ERROR: Drive %c: could not be found. Perhaps your hard disk needs to be partitioned first. Please create at least one primary partition on your hard disk, so SvarDOS can be installed on it. Note, that SvarDOS requires at least %d MiB of available disk space.\n\nYou can use the FDISK partitioning tool for creating the required partition manually, or you can let the installer partitioning your disk automatically. You can also abort the installation to use any other partition manager of your choice.
3.0:FEL: Enhet %c: kunde inte hittas. Kanske din h�rddisk beh�ver partitioneras f�rst. V�nligen skapa minst en prim�r partition p� din h�rddisk, s� SvarDOS kan installeras p� den. N.B. att SvarDOS beh�ver minst %d MiB ledigt diskutrymme.\n\nDu kan anv�nda FDISK-partitioneringsverktyget f�r att skapa den n�dv�ndiga partitionen manuellt, eller s� kan du l�ta installationsprogrammet partitioner din disk automatiskt. Du kan ocks� avbryta installationen f�r att anv�nda en annan valfri partitionsmanager.
#3.1:Your computer will reboot now.
3.1:Din dator kommer att boota om nu.
#3.2:ERROR: Drive %c: is a removable device. Installation aborted.
3.2:FEL: Enhet %c: �r ett removable device. Installationen avbryts.
#3.3:ERROR: Drive %c: seems to be unformated. Do you wish to format it?
3.3:FEL: Enhet %c: verkar vara oformaterad.
#3.4:ERROR: Drive %c: is not big enough! SvarDOS requires a disk of at least %d MiB.
3.4:FEL: Enhet %c: �r inte tillr�ckligt stor! SvarDOS beh�ver en disk som �r minst %d MiB.
#3.5:ERROR: Drive %c: is not empty. SvarDOS must be installed on an empty disk.\n\nYou can format the disk now, to make it empty. Note however, that this will ERASE ALL CURRENT DATA on your disk.
3.5:FEL: Enhet %c: �r inte tom. SvarDOS m�ste installeras p� en tom disk.\n\nDu kan formatera disken nu, f�r att t�mma den. N.B. detta kommer att RADERA ALLT NUVARANDE DATA p� din disk.
#3.6:The installation of SvarDOS to %c: is about to begin.
3.6:Installationen av SvarDOS till %c: ska just b�rja.

### PACKAGES INSTALLATION ###
### PAKETINSTALLATION ###
# example: "Installing package 4/50: FDISK"
# exempel: "Installerar paketet 4/50: FDISK"
#4.0:Installing package %d/%d: %s
4.0:Installerar paketet %d/%d: %s

### END SCREEN ###
### AVSLUTNINGSSKÄRM ###
#(5.0:SvarDOS installation is over. Your computer will reboot now.\nPlease remove the installation disk from your drive.)
#5.0:Your computer will reboot now.\nPlease make sure to remove the installation media.
5.0:Din dator kommer att reboota nu.\nV�nligen se till att ta bort installationsmediet.
#5.1:SvarDOS installation is over. Please restart your computer now.
5.1:SvarDOS-installationen �r klar. Please restart your computer now.

### LOG IN WELCOME TEXT ONCE SYSTEM IS INSTALLED ###
### LOGINV�LKOMSTTEXT N�R SYSTEMET �R INSTALLERAT ###
#6.0:Welcome to SvarDOS! Type 'HELP' if you need help.
6.0:V�lkommen till SvarDOS! Skriv 'HELP' om du beh�ver hj�lp.
